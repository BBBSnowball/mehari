../../../../../float_helpers.vhd