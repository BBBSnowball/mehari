../reconos/reconos/pcores/reconos_test_v3_01_a/hdl/vhdl/test_helpers.vhd