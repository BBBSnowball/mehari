../../../../../dummy_mod.vhd