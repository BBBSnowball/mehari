../../../../../float_neg.vhd