../../../../../double_type.vhd