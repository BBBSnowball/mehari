../../../../../float_sin.vhd