../../../../../single_pendulum.vhd