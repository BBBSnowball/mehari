../../../../../float_cos.vhd