../../../../../float_pkg_c_min.vhd